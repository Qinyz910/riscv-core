// Copyright (c) 2024
// SPDX-License-Identifier: Apache-2.0

`timescale 1ns/1ps

import rv32i_wb_pkg::*;

module rv32i_wb_data_adapter #(
  parameter int unsigned ADDR_WIDTH = WB_ADDR_WIDTH,
  parameter int unsigned DATA_WIDTH = WB_DATA_WIDTH
) (
  input  logic                     clk_i,
  input  logic                     rst_ni,

  // Pipeline side (MEM stage)
  input  logic                     req_i,
  input  logic                     we_i,
  input  logic [DATA_WIDTH/8-1:0]  be_i,
  input  logic [ADDR_WIDTH-1:0]    addr_i,
  input  logic [DATA_WIDTH-1:0]    wdata_i,
  output logic                     gnt_o,
  output logic                     rsp_valid_o,
  output logic [DATA_WIDTH-1:0]    rsp_rdata_o,
  output logic                     rsp_err_o,
  output logic                     store_complete_o,
  output logic                     store_err_o,

  // Wishbone master interface
  output logic                     wb_cyc_o,
  output logic                     wb_stb_o,
  output logic                     wb_we_o,
  output logic [DATA_WIDTH/8-1:0]  wb_sel_o,
  output logic [ADDR_WIDTH-1:0]    wb_adr_o,
  output logic [DATA_WIDTH-1:0]    wb_dat_o,
  input  logic [DATA_WIDTH-1:0]    wb_dat_i,
  input  logic                     wb_ack_i,
  input  logic                     wb_err_i,
  input  logic                     wb_stall_i
);

  logic                       pending_q;
  logic                       is_store_q;
  logic [ADDR_WIDTH-1:0]      addr_q;
  logic [DATA_WIDTH-1:0]      wdata_q;
  logic [DATA_WIDTH/8-1:0]    sel_q;

  logic                       rsp_valid_q;
  logic [DATA_WIDTH-1:0]      rsp_rdata_q;
  logic                       rsp_err_q;
  logic                       store_complete_q;
  logic                       store_err_q;

  logic accept_req;
  logic complete_transfer;

  assign accept_req        = (!pending_q) && req_i && !wb_stall_i;
  assign complete_transfer = pending_q && (wb_ack_i || wb_err_i);

  assign gnt_o             = accept_req;

  // Wishbone command outputs
  assign wb_cyc_o  = pending_q;
  assign wb_stb_o  = pending_q;
  assign wb_we_o   = is_store_q;
  assign wb_sel_o  = sel_q;
  assign wb_adr_o  = addr_q;
  assign wb_dat_o  = wdata_q;

  // Response outputs
  assign rsp_valid_o       = rsp_valid_q;
  assign rsp_rdata_o       = rsp_rdata_q;
  assign rsp_err_o         = rsp_err_q;
  assign store_complete_o  = store_complete_q;
  assign store_err_o       = store_err_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      pending_q          <= 1'b0;
      is_store_q         <= 1'b0;
      addr_q             <= '0;
      wdata_q            <= '0;
      sel_q              <= '0;
      rsp_valid_q        <= 1'b0;
      rsp_rdata_q        <= '0;
      rsp_err_q          <= 1'b0;
      store_complete_q   <= 1'b0;
      store_err_q        <= 1'b0;
    end else begin
      rsp_valid_q      <= 1'b0;
      store_complete_q <= 1'b0;
      store_err_q      <= 1'b0;

      if (accept_req) begin
        pending_q  <= 1'b1;
        is_store_q <= we_i;
        addr_q     <= addr_i;
        wdata_q    <= wdata_i;
        sel_q      <= we_i ? be_i : {DATA_WIDTH/8{1'b1}};
        rsp_err_q  <= 1'b0;
      end else if (complete_transfer) begin
        pending_q <= 1'b0;
        if (is_store_q) begin
          store_complete_q <= 1'b1;
          store_err_q      <= wb_err_i;
          rsp_err_q        <= 1'b0;
        end else begin
          rsp_valid_q <= 1'b1;
          rsp_err_q   <= wb_err_i;
          rsp_rdata_q <= wb_dat_i;
        end
      end
    end
  end

  // ---------------------------------------------------------------------------
  // Assertions
  // ---------------------------------------------------------------------------

  property p_no_overlap;
    @(posedge clk_i) disable iff (!rst_ni)
      pending_q |-> !accept_req;
  endproperty
  assert property (p_no_overlap)
    else $fatal(1, "[rv32i_wb_data_adapter] Overlapping data requests detected");

  property p_ack_only_when_pending;
    @(posedge clk_i) disable iff (!rst_ni)
      (wb_ack_i || wb_err_i) |-> pending_q;
  endproperty
  assert property (p_ack_only_when_pending)
    else $fatal(1, "[rv32i_wb_data_adapter] Response observed without an active transaction");

endmodule : rv32i_wb_data_adapter
